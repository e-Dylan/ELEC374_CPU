`timescale 1ns / 1ps

module and32(
	input wire [31:0] Ra,
	input wire [31:0] Rb,
	output wire [31:0] Rz
	);
	
	always @(*)
		assign RZ = Ra & Rb
endmodule

	