`timescale 1ns / 1ps

module negate32(
	input wire [31:0] Ra,
	output wire [31:0] Rz
	);
	
	wire [31:0] temp; 
	wire cout;
	not32 not_op(.Ra(Ra),.Rz(temp));
	add_32_bit add_op(.Ra(temp), .Rb(32'd1), .cin(1'd0),.sum(Rz), .cout(cout));
	
endmodule